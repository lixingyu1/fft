module rom_crtl (
    input                   clk,
    input                   rstn
);




endmodule //rom_crtl